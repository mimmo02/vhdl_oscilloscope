library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity test_signal is
    port (  clk_148_5_MHz   : in std_logic;
            reset           : in std_logic;
            
            next_sample : in std_logic;
            address     : out std_logic_vector(9 downto 0);
            data        : out std_logic_vector(19 downto 0));
end entity test_signal;

architecture platform_independent of test_signal is

    signal s_address : unsigned(9 downto 0);

begin

    address <= std_logic_vector(s_address);

    addr : process (clk_148_5_MHz, reset) is
    begin
        if reset = '1' THEN
            s_address <= ((others => '0'));
        elsif rising_edge(clk_148_5_MHz) THEN
            if next_sample = '1' then    
                s_address <= s_address + 1;
            end if;
        end if; 
    end process addr;

    rom : process (s_address) is
    begin
        case s_address is
            when "0000000000" => data <= "10000000001111111111";
            when "0000000001" => data <= "10000000111111110101";
            when "0000000010" => data <= "10000001101111010111";
            when "0000000011" => data <= "10000010011110100111";
            when "0000000100" => data <= "10000011001101100111";
            when "0000000101" => data <= "10000011111100011001";
            when "0000000110" => data <= "10000100101011000001";
            when "0000000111" => data <= "10000101011001100010";
            when "0000001000" => data <= "10000110011000000000";
            when "0000001001" => data <= "10000111000110011101";
            when "0000001010" => data <= "10000111110100111111";
            when "0000001011" => data <= "10001000100011101001";
            when "0000001100" => data <= "10001001010010011110";
            when "0000001101" => data <= "10001010000001100000";
            when "0000001110" => data <= "10001010110000110011";
            when "0000001111" => data <= "10001011110000011000";
            when "0000010000" => data <= "10001100100000001111";
            when "0000010001" => data <= "10001101010000011010";
            when "0000010010" => data <= "10001110000000110111";
            when "0000010011" => data <= "10001110110001100101";
            when "0000010100" => data <= "10001111100010100011";
            when "0000010101" => data <= "10010000010011101110";
            when "0000010110" => data <= "10010001000101000100";
            when "0000010111" => data <= "10010010000110100000";
            when "0000011000" => data <= "10010010110111111111";
            when "0000011001" => data <= "10010011101001011111";
            when "0000011010" => data <= "10010100011010111010";
            when "0000011011" => data <= "10010101001100001101";
            when "0000011100" => data <= "10010101111101010110";
            when "0000011101" => data <= "10010110101110010010";
            when "0000011110" => data <= "10010111011110111110";
            when "0000011111" => data <= "10011000001111011000";
            when "0000100000" => data <= "10011000111111100000";
            when "0000100001" => data <= "10011001101111010110";
            when "0000100010" => data <= "10011010101110111010";
            when "0000100011" => data <= "10011011011110001101";
            when "0000100100" => data <= "10011100001101010001";
            when "0000100101" => data <= "10011100111100001000";
            when "0000100110" => data <= "10011101101010110101";
            when "0000100111" => data <= "10011110011001011100";
            when "0000101000" => data <= "10011111001000000000";
            when "0000101001" => data <= "10011111110110100011";
            when "0000101010" => data <= "10100000100101001011";
            when "0000101011" => data <= "10100001010011111010";
            when "0000101100" => data <= "10100010000010110011";
            when "0000101101" => data <= "10100010110001111010";
            when "0000101110" => data <= "10100011100001001111";
            when "0000101111" => data <= "10100100010000110101";
            when "0000110000" => data <= "10100101000000101101";
            when "0000110001" => data <= "10100101110000110111";
            when "0000110010" => data <= "10100110100001010010";
            when "0000110011" => data <= "10100111010001111110";
            when "0000110100" => data <= "10101000000010111000";
            when "0000110101" => data <= "10101000110011111111";
            when "0000110110" => data <= "10101001100101001111";
            when "0000110111" => data <= "10101010010110100110";
            when "0000111000" => data <= "10101011000111111111";
            when "0000111001" => data <= "10101011111001011001";
            when "0000111010" => data <= "10101100101010101110";
            when "0000111011" => data <= "10101101011011111101";
            when "0000111100" => data <= "10101110001101000010";
            when "0000111101" => data <= "10101110111101111001";
            when "0000111110" => data <= "10101111101110100011";
            when "0000111111" => data <= "10110000011110111100";
            when "0001000000" => data <= "10110000111111000011";
            when "0001000001" => data <= "10110001101110111010";
            when "0001000010" => data <= "10110010011110011111";
            when "0001000011" => data <= "10110011001101110101";
            when "0001000100" => data <= "10110011111100111101";
            when "0001000101" => data <= "10110100101011111000";
            when "0001000110" => data <= "10110101011010101010";
            when "0001000111" => data <= "10110110001001010110";
            when "0001001000" => data <= "10110110101000000000";
            when "0001001001" => data <= "10110111010110101001";
            when "0001001010" => data <= "10111000000101010110";
            when "0001001011" => data <= "10111000110100001010";
            when "0001001100" => data <= "10111001100011000111";
            when "0001001101" => data <= "10111010010010010001";
            when "0001001110" => data <= "10111010110001101001";
            when "0001001111" => data <= "10111011100001010001";
            when "0001010000" => data <= "10111100010001001010";
            when "0001010001" => data <= "10111101000001010011";
            when "0001010010" => data <= "10111101100001101100";
            when "0001010011" => data <= "10111110010010010101";
            when "0001010100" => data <= "10111111000011001100";
            when "0001010101" => data <= "10111111110100001111";
            when "0001010110" => data <= "11000000010101011010";
            when "0001010111" => data <= "11000001000110101011";
            when "0001011000" => data <= "11000001110111111111";
            when "0001011001" => data <= "11000010011001010011";
            when "0001011010" => data <= "11000011001010100100";
            when "0001011011" => data <= "11000011111011101110";
            when "0001011100" => data <= "11000100011100101110";
            when "0001011101" => data <= "11000101001101100011";
            when "0001011110" => data <= "11000101111110001001";
            when "0001011111" => data <= "11000110011110100001";
            when "0001100000" => data <= "11000111001110101000";
            when "0001100001" => data <= "11000111111110011111";
            when "0001100010" => data <= "11001000011110000110";
            when "0001100011" => data <= "11001001001101011110";
            when "0001100100" => data <= "11001001101100101001";
            when "0001100101" => data <= "11001010011011101001";
            when "0001100110" => data <= "11001010111010100000";
            when "0001100111" => data <= "11001011101001010001";
            when "0001101000" => data <= "11001100001000000000";
            when "0001101001" => data <= "11001100110110101110";
            when "0001101010" => data <= "11001101100101100000";
            when "0001101011" => data <= "11001110000100011001";
            when "0001101100" => data <= "11001110100011011010";
            when "0001101101" => data <= "11001111010010100111";
            when "0001101110" => data <= "11001111110010000010";
            when "0001101111" => data <= "11010000100001101011";
            when "0001110000" => data <= "11010001000001100100";
            when "0001110001" => data <= "11010001110001101101";
            when "0001110010" => data <= "11010010010010000101";
            when "0001110011" => data <= "11010011000010101011";
            when "0001110100" => data <= "11010011100011011111";
            when "0001110101" => data <= "11010100000100011101";
            when "0001110110" => data <= "11010100110101100100";
            when "0001110111" => data <= "11010101010110110000";
            when "0001111000" => data <= "11010101110111111111";
            when "0001111001" => data <= "11010110101001001110";
            when "0001111010" => data <= "11010111001010011010";
            when "0001111011" => data <= "11010111101011011111";
            when "0001111100" => data <= "11011000011100011100";
            when "0001111101" => data <= "11011000111101001101";
            when "0001111110" => data <= "11011001011101110001";
            when "0001111111" => data <= "11011001111110000111";
            when "0010000000" => data <= "11011010101110001110";
            when "0010000001" => data <= "11011011001110000110";
            when "0010000010" => data <= "11011011101101101110";
            when "0010000011" => data <= "11011100001101001001";
            when "0010000100" => data <= "11011100101100010111";
            when "0010000101" => data <= "11011101001011011011";
            when "0010000110" => data <= "11011101111010010110";
            when "0010000111" => data <= "11011110011001001100";
            when "0010001000" => data <= "11011110111000000000";
            when "0010001001" => data <= "11011111010110110011";
            when "0010001010" => data <= "11011111110101101010";
            when "0010001011" => data <= "11100000010100100111";
            when "0010001100" => data <= "11100000110011101100";
            when "0010001101" => data <= "11100001010010111100";
            when "0010001110" => data <= "11100001110010011001";
            when "0010001111" => data <= "11100010010010000100";
            when "0010010000" => data <= "11100010110001111101";
            when "0010010001" => data <= "11100011010010000101";
            when "0010010010" => data <= "11100011110010011100";
            when "0010010011" => data <= "11100100010011000000";
            when "0010010100" => data <= "11100100110011110000";
            when "0010010101" => data <= "11100101010100101011";
            when "0010010110" => data <= "11100101110101101101";
            when "0010010111" => data <= "11100110010110110101";
            when "0010011000" => data <= "11100110110111111111";
            when "0010011001" => data <= "11100111011001001010";
            when "0010011010" => data <= "11100111101010010001";
            when "0010011011" => data <= "11101000001011010010";
            when "0010011100" => data <= "11101000101100001010";
            when "0010011101" => data <= "11101001001100111001";
            when "0010011110" => data <= "11101001101101011011";
            when "0010011111" => data <= "11101001111101110000";
            when "0010100000" => data <= "11101010011101110110";
            when "0010100001" => data <= "11101010111101101110";
            when "0010100010" => data <= "11101011011101011000";
            when "0010100011" => data <= "11101011101100110101";
            when "0010100100" => data <= "11101100001100000110";
            when "0010100101" => data <= "11101100101011001110";
            when "0010100110" => data <= "11101100111010001101";
            when "0010100111" => data <= "11101101011001001000";
            when "0010101000" => data <= "11101101111000000000";
            when "0010101001" => data <= "11101110000110111000";
            when "0010101010" => data <= "11101110100101110011";
            when "0010101011" => data <= "11101110110100110100";
            when "0010101100" => data <= "11101111010011111101";
            when "0010101101" => data <= "11101111110011010000";
            when "0010101110" => data <= "11110000000010101111";
            when "0010101111" => data <= "11110000100010011011";
            when "0010110000" => data <= "11110000110010010100";
            when "0010110001" => data <= "11110001010010011100";
            when "0010110010" => data <= "11110001100010110001";
            when "0010110011" => data <= "11110001110011010011";
            when "0010110100" => data <= "11110010010100000001";
            when "0010110101" => data <= "11110010100100111000";
            when "0010110110" => data <= "11110011000101110110";
            when "0010110111" => data <= "11110011010110111010";
            when "0010111000" => data <= "11110011100111111111";
            when "0010111001" => data <= "11110100001001000101";
            when "0010111010" => data <= "11110100011010001000";
            when "0010111011" => data <= "11110100101011000101";
            when "0010111100" => data <= "11110101001011111010";
            when "0010111101" => data <= "11110101011100100110";
            when "0010111110" => data <= "11110101101101000110";
            when "0010111111" => data <= "11110101111101011001";
            when "0011000000" => data <= "11110110011101011111";
            when "0011000001" => data <= "11110110101101011000";
            when "0011000010" => data <= "11110110111101000011";
            when "0011000011" => data <= "11110111001100100010";
            when "0011000100" => data <= "11110111011011110110";
            when "0011000101" => data <= "11110111101011000001";
            when "0011000110" => data <= "11110111111010000101";
            when "0011000111" => data <= "11111000011001000011";
            when "0011001000" => data <= "11111000101000000000";
            when "0011001001" => data <= "11111000110110111100";
            when "0011001010" => data <= "11111001000101111011";
            when "0011001011" => data <= "11111001010101000000";
            when "0011001100" => data <= "11111001100100001100";
            when "0011001101" => data <= "11111001110011100010";
            when "0011001110" => data <= "11111010000011000011";
            when "0011001111" => data <= "11111010010010110000";
            when "0011010000" => data <= "11111010010010101010";
            when "0011010001" => data <= "11111010100010110010";
            when "0011010010" => data <= "11111010110011000110";
            when "0011010011" => data <= "11111011000011100110";
            when "0011010100" => data <= "11111011010100010000";
            when "0011010101" => data <= "11111011100101000100";
            when "0011010110" => data <= "11111011110101111111";
            when "0011010111" => data <= "11111011110110111110";
            when "0011011000" => data <= "11111100000111111111";
            when "0011011001" => data <= "11111100011001000001";
            when "0011011010" => data <= "11111100101001111111";
            when "0011011011" => data <= "11111100101010111001";
            when "0011011100" => data <= "11111100111011101011";
            when "0011011101" => data <= "11111101001100010100";
            when "0011011110" => data <= "11111101001100110010";
            when "0011011111" => data <= "11111101011101000100";
            when "0011100000" => data <= "11111101101101001010";
            when "0011100001" => data <= "11111101101101000011";
            when "0011100010" => data <= "11111101111100110000";
            when "0011100011" => data <= "11111101111100010001";
            when "0011100100" => data <= "11111110001011100111";
            when "0011100101" => data <= "11111110001010110101";
            when "0011100110" => data <= "11111110011001111101";
            when "0011100111" => data <= "11111110011000111111";
            when "0011101000" => data <= "11111110101000000000";
            when "0011101001" => data <= "11111110100111000000";
            when "0011101010" => data <= "11111110110110000011";
            when "0011101011" => data <= "11111110110101001100";
            when "0011101100" => data <= "11111111000100011011";
            when "0011101101" => data <= "11111111000011110100";
            when "0011101110" => data <= "11111111000011010110";
            when "0011101111" => data <= "11111111010011000101";
            when "0011110000" => data <= "11111111010010111111";
            when "0011110001" => data <= "11111111010011000110";
            when "0011110010" => data <= "11111111100011011001";
            when "0011110011" => data <= "11111111100011110111";
            when "0011110100" => data <= "11111111100100011111";
            when "0011110101" => data <= "11111111100101001111";
            when "0011110110" => data <= "11111111110110000110";
            when "0011110111" => data <= "11111111110111000010";
            when "0011111000" => data <= "11111111110111111111";
            when "0011111001" => data <= "11111111111000111101";
            when "0011111010" => data <= "11111111111001111000";
            when "0011111011" => data <= "11111111111010101110";
            when "0011111100" => data <= "11111111111011011101";
            when "0011111101" => data <= "11111111111100000011";
            when "0011111110" => data <= "11111111111100100000";
            when "0011111111" => data <= "11111111111100110001";
            when "0100000000" => data <= "11111111111100110110";
            when "0100000001" => data <= "11111111111100101111";
            when "0100000010" => data <= "11111111111100011101";
            when "0100000011" => data <= "11111111111100000000";
            when "0100000100" => data <= "11111111111011011001";
            when "0100000101" => data <= "11111111111010101010";
            when "0100000110" => data <= "11111111111001110101";
            when "0100000111" => data <= "11111111111000111011";
            when "0100001000" => data <= "11111111111000000000";
            when "0100001001" => data <= "11111111110111000100";
            when "0100001010" => data <= "11111111110110001011";
            when "0100001011" => data <= "11111111100101010111";
            when "0100001100" => data <= "11111111100100101001";
            when "0100001101" => data <= "11111111100100000100";
            when "0100001110" => data <= "11111111100011101000";
            when "0100001111" => data <= "11111111010011011000";
            when "0100010000" => data <= "11111111010011010011";
            when "0100010001" => data <= "11111111010011011001";
            when "0100010010" => data <= "11111111000011101011";
            when "0100010011" => data <= "11111111000100000111";
            when "0100010100" => data <= "11111111000100101100";
            when "0100010101" => data <= "11111110110101011010";
            when "0100010110" => data <= "11111110110110001110";
            when "0100010111" => data <= "11111110100111000110";
            when "0100011000" => data <= "11111110100111111111";
            when "0100011001" => data <= "11111110011000111001";
            when "0100011010" => data <= "11111110011001110000";
            when "0100011011" => data <= "11111110001010100011";
            when "0100011100" => data <= "11111110001011001111";
            when "0100011101" => data <= "11111101111011110011";
            when "0100011110" => data <= "11111101111100001110";
            when "0100011111" => data <= "11111101101100011110";
            when "0100100000" => data <= "11111101101100100011";
            when "0100100001" => data <= "11111101011100011101";
            when "0100100010" => data <= "11111101001100001100";
            when "0100100011" => data <= "11111101001011110001";
            when "0100100100" => data <= "11111100111011001100";
            when "0100100101" => data <= "11111100101010100000";
            when "0100100110" => data <= "11111100101001101110";
            when "0100100111" => data <= "11111100011000111000";
            when "0100101000" => data <= "11111100001000000000";
            when "0100101001" => data <= "11111011110111001000";
            when "0100101010" => data <= "11111011110110010010";
            when "0100101011" => data <= "11111011100101100001";
            when "0100101100" => data <= "11111011010100110110";
            when "0100101101" => data <= "11111011000100010011";
            when "0100101110" => data <= "11111010110011111001";
            when "0100101111" => data <= "11111010100011101010";
            when "0100110000" => data <= "11111010010011100101";
            when "0100110001" => data <= "11111010010011101011";
            when "0100110010" => data <= "11111010000011111011";
            when "0100110011" => data <= "11111001110100010110";
            when "0100110100" => data <= "11111001100100111001";
            when "0100110101" => data <= "11111001010101100100";
            when "0100110110" => data <= "11111001000110010101";
            when "0100110111" => data <= "11111000110111001001";
            when "0100111000" => data <= "11111000100111111111";
            when "0100111001" => data <= "11111000011000110110";
            when "0100111010" => data <= "11110111111001101010";
            when "0100111011" => data <= "11110111101010011001";
            when "0100111100" => data <= "11110111011011000011";
            when "0100111101" => data <= "11110111001011100101";
            when "0100111110" => data <= "11110110111011111110";
            when "0100111111" => data <= "11110110101100001101";
            when "0101000000" => data <= "11110110011100010010";
            when "0101000001" => data <= "11110101111100001100";
            when "0101000010" => data <= "11110101101011111100";
            when "0101000011" => data <= "11110101011011100010";
            when "0101000100" => data <= "11110101001011000000";
            when "0101000101" => data <= "11110100101010010110";
            when "0101000110" => data <= "11110100011001100111";
            when "0101000111" => data <= "11110100001000110100";
            when "0101001000" => data <= "11110011101000000000";
            when "0101001001" => data <= "11110011010111001011";
            when "0101001010" => data <= "11110011000110011001";
            when "0101001011" => data <= "11110010100101101010";
            when "0101001100" => data <= "11110010010101000010";
            when "0101001101" => data <= "11110001110100100001";
            when "0101001110" => data <= "11110001100100001001";
            when "0101001111" => data <= "11110001010011111010";
            when "0101010000" => data <= "11110000110011110110";
            when "0101010001" => data <= "11110000100011111011";
            when "0101010010" => data <= "11110000000100001011";
            when "0101010011" => data <= "11101111110100100100";
            when "0101010100" => data <= "11101111010101000101";
            when "0101010101" => data <= "11101110110101101101";
            when "0101010110" => data <= "11101110100110011011";
            when "0101010111" => data <= "11101110000111001100";
            when "0101011000" => data <= "11101101110111111111";
            when "0101011001" => data <= "11101101011000110010";
            when "0101011010" => data <= "11101100111001100011";
            when "0101011011" => data <= "11101100101010010000";
            when "0101011100" => data <= "11101100001010110111";
            when "0101011101" => data <= "11101011101011010111";
            when "0101011110" => data <= "11101011011011101110";
            when "0101011111" => data <= "11101010111011111100";
            when "0101100000" => data <= "11101010011100000001";
            when "0101100001" => data <= "11101001111011111100";
            when "0101100010" => data <= "11101001101011101100";
            when "0101100011" => data <= "11101001001011010100";
            when "0101100100" => data <= "11101000101010110100";
            when "0101100101" => data <= "11101000001010001101";
            when "0101100110" => data <= "11100111101001100001";
            when "0101100111" => data <= "11100111011000110001";
            when "0101101000" => data <= "11100110111000000000";
            when "0101101001" => data <= "11100110010111001110";
            when "0101101010" => data <= "11100101110110011111";
            when "0101101011" => data <= "11100101010101110100";
            when "0101101100" => data <= "11100100110101001110";
            when "0101101101" => data <= "11100100010100101111";
            when "0101101110" => data <= "11100011110100011000";
            when "0101101111" => data <= "11100011010100001010";
            when "0101110000" => data <= "11100010110100000110";
            when "0101110001" => data <= "11100010010100001011";
            when "0101110010" => data <= "11100001110100011010";
            when "0101110011" => data <= "11100001010100110001";
            when "0101110100" => data <= "11100000110101010000";
            when "0101110101" => data <= "11100000010101110110";
            when "0101110110" => data <= "11011111110110100001";
            when "0101110111" => data <= "11011111010111001111";
            when "0101111000" => data <= "11011110110111111111";
            when "0101111001" => data <= "11011110011000101111";
            when "0101111010" => data <= "11011101111001011101";
            when "0101111011" => data <= "11011101001010000111";
            when "0101111100" => data <= "11011100101010101100";
            when "0101111101" => data <= "11011100001011001010";
            when "0101111110" => data <= "11011011101011100000";
            when "0101111111" => data <= "11011011001011101101";
            when "0110000000" => data <= "11011010101011110001";
            when "0110000001" => data <= "11011001111011101100";
            when "0110000010" => data <= "11011001011011011110";
            when "0110000011" => data <= "11011000111011000111";
            when "0110000100" => data <= "11011000011010101001";
            when "0110000101" => data <= "11010111101010000101";
            when "0110000110" => data <= "11010111001001011011";
            when "0110000111" => data <= "11010110101000101110";
            when "0110001000" => data <= "11010101111000000000";
            when "0110001001" => data <= "11010101010111010001";
            when "0110001010" => data <= "11010100110110100101";
            when "0110001011" => data <= "11010100000101111100";
            when "0110001100" => data <= "11010011100101011000";
            when "0110001101" => data <= "11010011000100111011";
            when "0110001110" => data <= "11010010010100100110";
            when "0110001111" => data <= "11010001110100011001";
            when "0110010000" => data <= "11010001000100010101";
            when "0110010001" => data <= "11010000100100011010";
            when "0110010010" => data <= "11001111110100101000";
            when "0110010011" => data <= "11001111010100111110";
            when "0110010100" => data <= "11001110100101011011";
            when "0110010101" => data <= "11001110000101111111";
            when "0110010110" => data <= "11001101100110100111";
            when "0110010111" => data <= "11001100110111010010";
            when "0110011000" => data <= "11001100000111111111";
            when "0110011001" => data <= "11001011101000101100";
            when "0110011010" => data <= "11001010111001010111";
            when "0110011011" => data <= "11001010011001111111";
            when "0110011100" => data <= "11001001101010100001";
            when "0110011101" => data <= "11001001001010111110";
            when "0110011110" => data <= "11001000011011010010";
            when "0110011111" => data <= "11000111111011011111";
            when "0110100000" => data <= "11000111001011100011";
            when "0110100001" => data <= "11000110011011011110";
            when "0110100010" => data <= "11000101111011010001";
            when "0110100011" => data <= "11000101001010111011";
            when "0110100100" => data <= "11000100011010011111";
            when "0110100101" => data <= "11000011111001111100";
            when "0110100110" => data <= "11000011001001010101";
            when "0110100111" => data <= "11000010011000101011";
            when "0110101000" => data <= "11000001111000000000";
            when "0110101001" => data <= "11000001000111010100";
            when "0110101010" => data <= "11000000010110101010";
            when "0110101011" => data <= "10111111110110000100";
            when "0110101100" => data <= "10111111000101100011";
            when "0110101101" => data <= "10111110010101000111";
            when "0110101110" => data <= "10111101100100110011";
            when "0110101111" => data <= "10111101000100100111";
            when "0110110000" => data <= "10111100010100100011";
            when "0110110001" => data <= "10111011100100101000";
            when "0110110010" => data <= "10111010110100110101";
            when "0110110011" => data <= "10111010010101001001";
            when "0110110100" => data <= "10111001100101100101";
            when "0110110101" => data <= "10111000110110000110";
            when "0110110110" => data <= "10111000000110101100";
            when "0110110111" => data <= "10110111010111010101";
            when "0110111000" => data <= "10110110100111111111";
            when "0110111001" => data <= "10110110001000101010";
            when "0110111010" => data <= "10110101011001010010";
            when "0110111011" => data <= "10110100101001110111";
            when "0110111100" => data <= "10110011111010011000";
            when "0110111101" => data <= "10110011001010110010";
            when "0110111110" => data <= "10110010011011000101";
            when "0110111111" => data <= "10110001101011010001";
            when "0111000000" => data <= "10110000111011010101";
            when "0111000001" => data <= "10110000011011010000";
            when "0111000010" => data <= "10101111101011000100";
            when "0111000011" => data <= "10101110111010110000";
            when "0111000100" => data <= "10101110001010010101";
            when "0111000101" => data <= "10101101011001110101";
            when "0111000110" => data <= "10101100101001010000";
            when "0111000111" => data <= "10101011111000101001";
            when "0111001000" => data <= "10101011001000000000";
            when "0111001001" => data <= "10101010010111010111";
            when "0111001010" => data <= "10101001100110101111";
            when "0111001011" => data <= "10101000110110001011";
            when "0111001100" => data <= "10101000000101101100";
            when "0111001101" => data <= "10100111010101010010";
            when "0111001110" => data <= "10100110100101000000";
            when "0111001111" => data <= "10100101110100110100";
            when "0111010000" => data <= "10100101000100110001";
            when "0111010001" => data <= "10100100010100110101";
            when "0111010010" => data <= "10100011100101000001";
            when "0111010011" => data <= "10100010110101010101";
            when "0111010100" => data <= "10100010000101101110";
            when "0111010101" => data <= "10100001010110001110";
            when "0111010110" => data <= "10100000100110110001";
            when "0111010111" => data <= "10011111110111011000";
            when "0111011000" => data <= "10011111000111111111";
            when "0111011001" => data <= "10011110011000100111";
            when "0111011010" => data <= "10011101101001001101";
            when "0111011011" => data <= "10011100111001110000";
            when "0111011100" => data <= "10011100001010001110";
            when "0111011101" => data <= "10011011011010100111";
            when "0111011110" => data <= "10011010101010111001";
            when "0111011111" => data <= "10011001101011000101";
            when "0111100000" => data <= "10011000111011001000";
            when "0111100001" => data <= "10011000001011000100";
            when "0111100010" => data <= "10010111011010111000";
            when "0111100011" => data <= "10010110101010100101";
            when "0111100100" => data <= "10010101111010001100";
            when "0111100101" => data <= "10010101001001101110";
            when "0111100110" => data <= "10010100011001001011";
            when "0111100111" => data <= "10010011101000100110";
            when "0111101000" => data <= "10010010111000000000";
            when "0111101001" => data <= "10010010000111011001";
            when "0111101010" => data <= "10010001000110110100";
            when "0111101011" => data <= "10010000010110010010";
            when "0111101100" => data <= "10001111100101110101";
            when "0111101101" => data <= "10001110110101011101";
            when "0111101110" => data <= "10001110000101001011";
            when "0111101111" => data <= "10001101010101000001";
            when "0111110000" => data <= "10001100100100111101";
            when "0111110001" => data <= "10001011110101000001";
            when "0111110010" => data <= "10001010110101001101";
            when "0111110011" => data <= "10001010000101011111";
            when "0111110100" => data <= "10001001010101110111";
            when "0111110101" => data <= "10001000100110010101";
            when "0111110110" => data <= "10000111110110110110";
            when "0111110111" => data <= "10000111000111011010";
            when "0111111000" => data <= "10000110010111111111";
            when "0111111001" => data <= "10000101011000100101";
            when "0111111010" => data <= "10000100101001001000";
            when "0111111011" => data <= "10000011111001101001";
            when "0111111100" => data <= "10000011001010000110";
            when "0111111101" => data <= "10000010011010011101";
            when "0111111110" => data <= "10000001101010101110";
            when "0111111111" => data <= "10000000111010111001";
            when "1000000000" => data <= "10000000001010111100";
            when "1000000001" => data <= "01111111001010111000";
            when "1000000010" => data <= "01111110011010101101";
            when "1000000011" => data <= "01111101101010011011";
            when "1000000100" => data <= "01111100111010000100";
            when "1000000101" => data <= "01111100001001100111";
            when "1000000110" => data <= "01111011011001000111";
            when "1000000111" => data <= "01111010101000100100";
            when "1000001000" => data <= "01111001101000000000";
            when "1000001001" => data <= "01111000110111011011";
            when "1000001010" => data <= "01111000000110111001";
            when "1000001011" => data <= "01110111010110011001";
            when "1000001100" => data <= "01110110100101111101";
            when "1000001101" => data <= "01110101110101100111";
            when "1000001110" => data <= "01110101000101010110";
            when "1000001111" => data <= "01110100000101001100";
            when "1000010000" => data <= "01110011010101001001";
            when "1000010001" => data <= "01110010100101001101";
            when "1000010010" => data <= "01110001110101010111";
            when "1000010011" => data <= "01110001000101101001";
            when "1000010100" => data <= "01110000010101111111";
            when "1000010101" => data <= "01101111100110011011";
            when "1000010110" => data <= "01101110110110111010";
            when "1000010111" => data <= "01101101110111011100";
            when "1000011000" => data <= "01101101000111111111";
            when "1000011001" => data <= "01101100011000100010";
            when "1000011010" => data <= "01101011101001000100";
            when "1000011011" => data <= "01101010111001100011";
            when "1000011100" => data <= "01101010001001111110";
            when "1000011101" => data <= "01101001011010010011";
            when "1000011110" => data <= "01101000101010100100";
            when "1000011111" => data <= "01100111111010101101";
            when "1000100000" => data <= "01100111001010110000";
            when "1000100001" => data <= "01100110011010101101";
            when "1000100010" => data <= "01100101011010100010";
            when "1000100011" => data <= "01100100101010010010";
            when "1000100100" => data <= "01100011111001111100";
            when "1000100101" => data <= "01100011001001100001";
            when "1000100110" => data <= "01100010011001000010";
            when "1000100111" => data <= "01100001101000100010";
            when "1000101000" => data <= "01100000111000000000";
            when "1000101001" => data <= "01100000000111011110";
            when "1000101010" => data <= "01011111010110111101";
            when "1000101011" => data <= "01011110100110011111";
            when "1000101100" => data <= "01011101110110000101";
            when "1000101101" => data <= "01011101000101110000";
            when "1000101110" => data <= "01011100010101100000";
            when "1000101111" => data <= "01011011100101010111";
            when "1000110000" => data <= "01011010110101010100";
            when "1000110001" => data <= "01011010000101011000";
            when "1000110010" => data <= "01011001010101100010";
            when "1000110011" => data <= "01011000100101110010";
            when "1000110100" => data <= "01010111110110000111";
            when "1000110101" => data <= "01010111000110100001";
            when "1000110110" => data <= "01010110010110111111";
            when "1000110111" => data <= "01010101100111011110";
            when "1000111000" => data <= "01010100110111111111";
            when "1000111001" => data <= "01010100001000100000";
            when "1000111010" => data <= "01010011011001000000";
            when "1000111011" => data <= "01010010101001011101";
            when "1000111100" => data <= "01010001111001110110";
            when "1000111101" => data <= "01010001001010001011";
            when "1000111110" => data <= "01010000011010011010";
            when "1000111111" => data <= "01001111101010100011";
            when "1001000000" => data <= "01001111001010100110";
            when "1001000001" => data <= "01001110011010100010";
            when "1001000010" => data <= "01001101101010011000";
            when "1001000011" => data <= "01001100111010001001";
            when "1001000100" => data <= "01001100001001110100";
            when "1001000101" => data <= "01001011011001011011";
            when "1001000110" => data <= "01001010101000111110";
            when "1001000111" => data <= "01001001111000011111";
            when "1001001000" => data <= "01001001011000000000";
            when "1001001001" => data <= "01001000100111100000";
            when "1001001010" => data <= "01000111110111000001";
            when "1001001011" => data <= "01000111000110100101";
            when "1001001100" => data <= "01000110010110001101";
            when "1001001101" => data <= "01000101100101111001";
            when "1001001110" => data <= "01000101000101101010";
            when "1001001111" => data <= "01000100010101100001";
            when "1001010000" => data <= "01000011100101011110";
            when "1001010001" => data <= "01000010110101100010";
            when "1001010010" => data <= "01000010010101101011";
            when "1001010011" => data <= "01000001100101111010";
            when "1001010100" => data <= "01000000110110001110";
            when "1001010101" => data <= "01000000000110100111";
            when "1001010110" => data <= "00111111100111000011";
            when "1001010111" => data <= "00111110110111100000";
            when "1001011000" => data <= "00111110000111111111";
            when "1001011001" => data <= "00111101101000011110";
            when "1001011010" => data <= "00111100111000111100";
            when "1001011011" => data <= "00111100001001010111";
            when "1001011100" => data <= "00111011101001101111";
            when "1001011101" => data <= "00111010111010000010";
            when "1001011110" => data <= "00111010001010010000";
            when "1001011111" => data <= "00111001101010011001";
            when "1001100000" => data <= "00111000111010011100";
            when "1001100001" => data <= "00111000001010011000";
            when "1001100010" => data <= "00110111101010001111";
            when "1001100011" => data <= "00110110111010000001";
            when "1001100100" => data <= "00110110011001101101";
            when "1001100101" => data <= "00110101101001010101";
            when "1001100110" => data <= "00110101001000111011";
            when "1001100111" => data <= "00110100011000011110";
            when "1001101000" => data <= "00110011111000000000";
            when "1001101001" => data <= "00110011000111100010";
            when "1001101010" => data <= "00110010010111000101";
            when "1001101011" => data <= "00110001110110101011";
            when "1001101100" => data <= "00110001010110010100";
            when "1001101101" => data <= "00110000100110000001";
            when "1001101110" => data <= "00110000000101110011";
            when "1001101111" => data <= "00101111010101101011";
            when "1001110000" => data <= "00101110110101101000";
            when "1001110001" => data <= "00101110000101101011";
            when "1001110010" => data <= "00101101100101110100";
            when "1001110011" => data <= "00101100110110000010";
            when "1001110100" => data <= "00101100010110010101";
            when "1001110101" => data <= "00101011110110101100";
            when "1001110110" => data <= "00101011000111000110";
            when "1001110111" => data <= "00101010100111100010";
            when "1001111000" => data <= "00101010000111111111";
            when "1001111001" => data <= "00101001011000011101";
            when "1001111010" => data <= "00101000111000111000";
            when "1001111011" => data <= "00101000011001010010";
            when "1001111100" => data <= "00100111101001101000";
            when "1001111101" => data <= "00100111001001111010";
            when "1001111110" => data <= "00100110101010001000";
            when "1001111111" => data <= "00100110001010010000";
            when "1010000000" => data <= "00100101011010010010";
            when "1010000001" => data <= "00100100111010001111";
            when "1010000010" => data <= "00100100011010000110";
            when "1010000011" => data <= "00100011111001111001";
            when "1010000100" => data <= "00100011011001100110";
            when "1010000101" => data <= "00100010111001010000";
            when "1010000110" => data <= "00100010001000110111";
            when "1010000111" => data <= "00100001101000011100";
            when "1010001000" => data <= "00100001001000000000";
            when "1010001001" => data <= "00100000100111100011";
            when "1010001010" => data <= "00100000000111001000";
            when "1010001011" => data <= "00011111100110110000";
            when "1010001100" => data <= "00011111000110011010";
            when "1010001101" => data <= "00011110100110001001";
            when "1010001110" => data <= "00011110000101111100";
            when "1010001111" => data <= "00011101100101110100";
            when "1010010000" => data <= "00011101000101110001";
            when "1010010001" => data <= "00011100100101110100";
            when "1010010010" => data <= "00011100000101111101";
            when "1010010011" => data <= "00011011100110001010";
            when "1010010100" => data <= "00011011000110011100";
            when "1010010101" => data <= "00011010100110110001";
            when "1010010110" => data <= "00011010000111001010";
            when "1010010111" => data <= "00011001100111100100";
            when "1010011000" => data <= "00011001000111111111";
            when "1010011001" => data <= "00011000101000011011";
            when "1010011010" => data <= "00011000011000110101";
            when "1010011011" => data <= "00010111111001001101";
            when "1010011100" => data <= "00010111011001100010";
            when "1010011101" => data <= "00010110111001110011";
            when "1010011110" => data <= "00010110011001111111";
            when "1010011111" => data <= "00010110001010000111";
            when "1010100000" => data <= "00010101101010001001";
            when "1010100001" => data <= "00010101001010000110";
            when "1010100010" => data <= "00010100101001111110";
            when "1010100011" => data <= "00010100011001110001";
            when "1010100100" => data <= "00010011111001100000";
            when "1010100101" => data <= "00010011011001001011";
            when "1010100110" => data <= "00010011001000110100";
            when "1010100111" => data <= "00010010101000011010";
            when "1010101000" => data <= "00010010001000000000";
            when "1010101001" => data <= "00010001110111100101";
            when "1010101010" => data <= "00010001010111001100";
            when "1010101011" => data <= "00010001000110110101";
            when "1010101100" => data <= "00010000100110100000";
            when "1010101101" => data <= "00010000000110010000";
            when "1010101110" => data <= "00001111110110000100";
            when "1010101111" => data <= "00001111010101111100";
            when "1010110000" => data <= "00001111000101111010";
            when "1010110001" => data <= "00001110100101111101";
            when "1010110010" => data <= "00001110010110000101";
            when "1010110011" => data <= "00001110000110010001";
            when "1010110100" => data <= "00001101100110100010";
            when "1010110101" => data <= "00001101010110110110";
            when "1010110110" => data <= "00001100110111001101";
            when "1010110111" => data <= "00001100100111100110";
            when "1010111000" => data <= "00001100010111111111";
            when "1010111001" => data <= "00001011111000011001";
            when "1010111010" => data <= "00001011101000110010";
            when "1010111011" => data <= "00001011011001001000";
            when "1010111100" => data <= "00001010111001011100";
            when "1010111101" => data <= "00001010101001101100";
            when "1010111110" => data <= "00001010011001111000";
            when "1010111111" => data <= "00001010001001111111";
            when "1011000000" => data <= "00001001101010000001";
            when "1011000001" => data <= "00001001011001111110";
            when "1011000010" => data <= "00001001001001110111";
            when "1011000011" => data <= "00001000111001101011";
            when "1011000100" => data <= "00001000101001011010";
            when "1011000101" => data <= "00001000011001000111";
            when "1011000110" => data <= "00001000001000110000";
            when "1011000111" => data <= "00000111101000011000";
            when "1011001000" => data <= "00000111011000000000";
            when "1011001001" => data <= "00000111000111100111";
            when "1011001010" => data <= "00000110110111001111";
            when "1011001011" => data <= "00000110100110111001";
            when "1011001100" => data <= "00000110010110100110";
            when "1011001101" => data <= "00000110000110010111";
            when "1011001110" => data <= "00000101110110001011";
            when "1011001111" => data <= "00000101100110000100";
            when "1011010000" => data <= "00000101100110000010";
            when "1011010001" => data <= "00000101010110000101";
            when "1011010010" => data <= "00000101000110001100";
            when "1011010011" => data <= "00000100110110011000";
            when "1011010100" => data <= "00000100100110100111";
            when "1011010101" => data <= "00000100010110111010";
            when "1011010110" => data <= "00000100000111010000";
            when "1011010111" => data <= "00000100000111100111";
            when "1011011000" => data <= "00000011110111111111";
            when "1011011001" => data <= "00000011101000011000";
            when "1011011010" => data <= "00000011011000101111";
            when "1011011011" => data <= "00000011011001000100";
            when "1011011100" => data <= "00000011001001010110";
            when "1011011101" => data <= "00000010111001100101";
            when "1011011110" => data <= "00000010111001110000";
            when "1011011111" => data <= "00000010101001110111";
            when "1011100000" => data <= "00000010011001111001";
            when "1011100001" => data <= "00000010011001110111";
            when "1011100010" => data <= "00000010001001101111";
            when "1011100011" => data <= "00000010001001100100";
            when "1011100100" => data <= "00000001111001010101";
            when "1011100101" => data <= "00000001111001000010";
            when "1011100110" => data <= "00000001101000101101";
            when "1011100111" => data <= "00000001101000010111";
            when "1011101000" => data <= "00000001011000000000";
            when "1011101001" => data <= "00000001010111101000";
            when "1011101010" => data <= "00000001000111010010";
            when "1011101011" => data <= "00000001000110111101";
            when "1011101100" => data <= "00000000110110101100";
            when "1011101101" => data <= "00000000110110011101";
            when "1011101110" => data <= "00000000110110010010";
            when "1011101111" => data <= "00000000100110001100";
            when "1011110000" => data <= "00000000100110001010";
            when "1011110001" => data <= "00000000100110001100";
            when "1011110010" => data <= "00000000010110010011";
            when "1011110011" => data <= "00000000010110011110";
            when "1011110100" => data <= "00000000010110101101";
            when "1011110101" => data <= "00000000010110111111";
            when "1011110110" => data <= "00000000000111010011";
            when "1011110111" => data <= "00000000000111101001";
            when "1011111000" => data <= "00000000000111111111";
            when "1011111001" => data <= "00000000001000010110";
            when "1011111010" => data <= "00000000001000101100";
            when "1011111011" => data <= "00000000001001000000";
            when "1011111100" => data <= "00000000001001010001";
            when "1011111101" => data <= "00000000001001011111";
            when "1011111110" => data <= "00000000001001101001";
            when "1011111111" => data <= "00000000001001110000";
            when "1100000000" => data <= "00000000001001110010";
            when "1100000001" => data <= "00000000001001101111";
            when "1100000010" => data <= "00000000001001101001";
            when "1100000011" => data <= "00000000001001011110";
            when "1100000100" => data <= "00000000001001010000";
            when "1100000101" => data <= "00000000001000111110";
            when "1100000110" => data <= "00000000001000101011";
            when "1100000111" => data <= "00000000001000010101";
            when "1100001000" => data <= "00000000001000000000";
            when "1100001001" => data <= "00000000000111101010";
            when "1100001010" => data <= "00000000000111010101";
            when "1100001011" => data <= "00000000010111000001";
            when "1100001100" => data <= "00000000010110110001";
            when "1100001101" => data <= "00000000010110100011";
            when "1100001110" => data <= "00000000010110011001";
            when "1100001111" => data <= "00000000100110010011";
            when "1100010000" => data <= "00000000100110010001";
            when "1100010001" => data <= "00000000100110010011";
            when "1100010010" => data <= "00000000110110011010";
            when "1100010011" => data <= "00000000110110100100";
            when "1100010100" => data <= "00000000110110110010";
            when "1100010101" => data <= "00000001000111000011";
            when "1100010110" => data <= "00000001000111010110";
            when "1100010111" => data <= "00000001010111101010";
            when "1100011000" => data <= "00000001010111111111";
            when "1100011001" => data <= "00000001101000010101";
            when "1100011010" => data <= "00000001101000101001";
            when "1100011011" => data <= "00000001111000111100";
            when "1100011100" => data <= "00000001111001001100";
            when "1100011101" => data <= "00000010001001011001";
            when "1100011110" => data <= "00000010001001100011";
            when "1100011111" => data <= "00000010011001101001";
            when "1100100000" => data <= "00000010011001101011";
            when "1100100001" => data <= "00000010101001101001";
            when "1100100010" => data <= "00000010111001100010";
            when "1100100011" => data <= "00000010111001011000";
            when "1100100100" => data <= "00000011001001001011";
            when "1100100101" => data <= "00000011011000111011";
            when "1100100110" => data <= "00000011011000101000";
            when "1100100111" => data <= "00000011101000010100";
            when "1100101000" => data <= "00000011111000000000";
            when "1100101001" => data <= "00000100000111101011";
            when "1100101010" => data <= "00000100000111010111";
            when "1100101011" => data <= "00000100010111000101";
            when "1100101100" => data <= "00000100100110110101";
            when "1100101101" => data <= "00000100110110101001";
            when "1100101110" => data <= "00000101000110011111";
            when "1100101111" => data <= "00000101010110011001";
            when "1100110000" => data <= "00000101100110010111";
            when "1100110001" => data <= "00000101100110011010";
            when "1100110010" => data <= "00000101110110100000";
            when "1100110011" => data <= "00000110000110101010";
            when "1100110100" => data <= "00000110010110110111";
            when "1100110101" => data <= "00000110100111000110";
            when "1100110110" => data <= "00000110110111011000";
            when "1100110111" => data <= "00000111000111101011";
            when "1100111000" => data <= "00000111010111111111";
            when "1100111001" => data <= "00000111101000010011";
            when "1100111010" => data <= "00001000001000100111";
            when "1100111011" => data <= "00001000011000111000";
            when "1100111100" => data <= "00001000101001000111";
            when "1100111101" => data <= "00001000111001010100";
            when "1100111110" => data <= "00001001001001011101";
            when "1100111111" => data <= "00001001011001100011";
            when "1101000000" => data <= "00001001101001100100";
            when "1101000001" => data <= "00001010001001100010";
            when "1101000010" => data <= "00001010011001011100";
            when "1101000011" => data <= "00001010101001010011";
            when "1101000100" => data <= "00001010111001000110";
            when "1101000101" => data <= "00001011011000110111";
            when "1101000110" => data <= "00001011101000100110";
            when "1101000111" => data <= "00001011111000010011";
            when "1101001000" => data <= "00001100011000000000";
            when "1101001001" => data <= "00001100100111101100";
            when "1101001010" => data <= "00001100110111011010";
            when "1101001011" => data <= "00001101010111001001";
            when "1101001100" => data <= "00001101100110111010";
            when "1101001101" => data <= "00001110000110101110";
            when "1101001110" => data <= "00001110010110100101";
            when "1101001111" => data <= "00001110100110011111";
            when "1101010000" => data <= "00001111000110011110";
            when "1101010001" => data <= "00001111010110100000";
            when "1101010010" => data <= "00001111110110100110";
            when "1101010011" => data <= "00010000000110101111";
            when "1101010100" => data <= "00010000100110111011";
            when "1101010101" => data <= "00010001000111001010";
            when "1101010110" => data <= "00010001010111011011";
            when "1101010111" => data <= "00010001110111101101";
            when "1101011000" => data <= "00010010000111111111";
            when "1101011001" => data <= "00010010101000010010";
            when "1101011010" => data <= "00010011001000100100";
            when "1101011011" => data <= "00010011011000110101";
            when "1101011100" => data <= "00010011111001000011";
            when "1101011101" => data <= "00010100011001001111";
            when "1101011110" => data <= "00010100101001010111";
            when "1101011111" => data <= "00010101001001011101";
            when "1101100000" => data <= "00010101101001011110";
            when "1101100001" => data <= "00010110001001011100";
            when "1101100010" => data <= "00010110011001010111";
            when "1101100011" => data <= "00010110111001001110";
            when "1101100100" => data <= "00010111011001000010";
            when "1101100101" => data <= "00010111111000110100";
            when "1101100110" => data <= "00011000011000100011";
            when "1101100111" => data <= "00011000101000010010";
            when "1101101000" => data <= "00011001001000000000";
            when "1101101001" => data <= "00011001100111101101";
            when "1101101010" => data <= "00011010000111011100";
            when "1101101011" => data <= "00011010100111001100";
            when "1101101100" => data <= "00011011000110111110";
            when "1101101101" => data <= "00011011100110110011";
            when "1101101110" => data <= "00011100000110101010";
            when "1101101111" => data <= "00011100100110100101";
            when "1101110000" => data <= "00011101000110100100";
            when "1101110001" => data <= "00011101100110100110";
            when "1101110010" => data <= "00011110000110101011";
            when "1101110011" => data <= "00011110100110110100";
            when "1101110100" => data <= "00011111000110111111";
            when "1101110101" => data <= "00011111100111001101";
            when "1101110110" => data <= "00100000000111011101";
            when "1101110111" => data <= "00100000100111101110";
            when "1101111000" => data <= "00100001000111111111";
            when "1101111001" => data <= "00100001101000010001";
            when "1101111010" => data <= "00100010001000100010";
            when "1101111011" => data <= "00100010111000110001";
            when "1101111100" => data <= "00100011011000111111";
            when "1101111101" => data <= "00100011111001001010";
            when "1101111110" => data <= "00100100011001010010";
            when "1101111111" => data <= "00100100111001010111";
            when "1110000000" => data <= "00100101011001011000";
            when "1110000001" => data <= "00100110001001010111";
            when "1110000010" => data <= "00100110101001010001";
            when "1110000011" => data <= "00100111001001001001";
            when "1110000100" => data <= "00100111101000111110";
            when "1110000101" => data <= "00101000011000110000";
            when "1110000110" => data <= "00101000111000100001";
            when "1110000111" => data <= "00101001011000010001";
            when "1110001000" => data <= "00101010001000000000";
            when "1110001001" => data <= "00101010100111101110";
            when "1110001010" => data <= "00101011000111011110";
            when "1110001011" => data <= "00101011110111001111";
            when "1110001100" => data <= "00101100010111000010";
            when "1110001101" => data <= "00101100110110110111";
            when "1110001110" => data <= "00101101100110110000";
            when "1110001111" => data <= "00101110000110101011";
            when "1110010000" => data <= "00101110110110101001";
            when "1110010001" => data <= "00101111010110101011";
            when "1110010010" => data <= "00110000000110110000";
            when "1110010011" => data <= "00110000100110111000";
            when "1110010100" => data <= "00110001010111000011";
            when "1110010101" => data <= "00110001110111010000";
            when "1110010110" => data <= "00110010010111011111";
            when "1110010111" => data <= "00110011000111101111";
            when "1110011000" => data <= "00110011110111111111";
            when "1110011001" => data <= "00110100011000010000";
            when "1110011010" => data <= "00110101001000100000";
            when "1110011011" => data <= "00110101101000101110";
            when "1110011100" => data <= "00110110011000111011";
            when "1110011101" => data <= "00110110111001000101";
            when "1110011110" => data <= "00110111101001001101";
            when "1110011111" => data <= "00111000001001010010";
            when "1110100000" => data <= "00111000111001010011";
            when "1110100001" => data <= "00111001101001010001";
            when "1110100010" => data <= "00111010001001001100";
            when "1110100011" => data <= "00111010111001000101";
            when "1110100100" => data <= "00111011101000111010";
            when "1110100101" => data <= "00111100001000101101";
            when "1110100110" => data <= "00111100111000011111";
            when "1110100111" => data <= "00111101101000010000";
            when "1110101000" => data <= "00111110001000000000";
            when "1110101001" => data <= "00111110110111101111";
            when "1110101010" => data <= "00111111100111100000";
            when "1110101011" => data <= "01000000000111010010";
            when "1110101100" => data <= "01000000110111000110";
            when "1110101101" => data <= "01000001100110111100";
            when "1110101110" => data <= "01000010010110110100";
            when "1110101111" => data <= "01000010110110110000";
            when "1110110000" => data <= "01000011100110101110";
            when "1110110001" => data <= "01000100010110110000";
            when "1110110010" => data <= "01000101000110110101";
            when "1110110011" => data <= "01000101100110111101";
            when "1110110100" => data <= "01000110010111000111";
            when "1110110101" => data <= "01000111000111010011";
            when "1110110110" => data <= "01000111110111100001";
            when "1110110111" => data <= "01001000100111110000";
            when "1110111000" => data <= "01001001010111111111";
            when "1110111001" => data <= "01001001111000001111";
            when "1110111010" => data <= "01001010101000011110";
            when "1110111011" => data <= "01001011011000101100";
            when "1110111100" => data <= "01001100001000110111";
            when "1110111101" => data <= "01001100111001000001";
            when "1110111110" => data <= "01001101101001001000";
            when "1110111111" => data <= "01001110011001001101";
            when "1111000000" => data <= "01001111001001001110";
            when "1111000001" => data <= "01001111101001001100";
            when "1111000010" => data <= "01010000011001001000";
            when "1111000011" => data <= "01010001001001000000";
            when "1111000100" => data <= "01010001111000110111";
            when "1111000101" => data <= "01010010101000101011";
            when "1111000110" => data <= "01010011011000011101";
            when "1111000111" => data <= "01010100001000001111";
            when "1111001000" => data <= "01010100111000000000";
            when "1111001001" => data <= "01010101100111110000";
            when "1111001010" => data <= "01010110010111100010";
            when "1111001011" => data <= "01010111000111010101";
            when "1111001100" => data <= "01010111110111001001";
            when "1111001101" => data <= "01011000100111000000";
            when "1111001110" => data <= "01011001010110111001";
            when "1111001111" => data <= "01011010000110110101";
            when "1111010000" => data <= "01011010110110110011";
            when "1111010001" => data <= "01011011100110110101";
            when "1111010010" => data <= "01011100010110111001";
            when "1111010011" => data <= "01011101000111000001";
            when "1111010100" => data <= "01011101110111001010";
            when "1111010101" => data <= "01011110100111010110";
            when "1111010110" => data <= "01011111010111100011";
            when "1111010111" => data <= "01100000000111110001";
            when "1111011000" => data <= "01100000110111111111";
            when "1111011001" => data <= "01100001101000001110";
            when "1111011010" => data <= "01100010011000011100";
            when "1111011011" => data <= "01100011001000101001";
            when "1111011100" => data <= "01100011111000110100";
            when "1111011101" => data <= "01100100101000111101";
            when "1111011110" => data <= "01100101011001000100";
            when "1111011111" => data <= "01100110011001001000";
            when "1111100000" => data <= "01100111001001001001";
            when "1111100001" => data <= "01100111111001001000";
            when "1111100010" => data <= "01101000101001000011";
            when "1111100011" => data <= "01101001011000111100";
            when "1111100100" => data <= "01101010001000110011";
            when "1111100101" => data <= "01101010111000101000";
            when "1111100110" => data <= "01101011101000011011";
            when "1111100111" => data <= "01101100011000001110";
            when "1111101000" => data <= "01101101001000000000";
            when "1111101001" => data <= "01101101110111110001";
            when "1111101010" => data <= "01101110110111100100";
            when "1111101011" => data <= "01101111100111010111";
            when "1111101100" => data <= "01110000010111001101";
            when "1111101101" => data <= "01110001000111000100";
            when "1111101110" => data <= "01110001110110111101";
            when "1111101111" => data <= "01110010100110111001";
            when "1111110000" => data <= "01110011010110111000";
            when "1111110001" => data <= "01110100000110111010";
            when "1111110010" => data <= "01110101000110111110";
            when "1111110011" => data <= "01110101110111000100";
            when "1111110100" => data <= "01110110100111001101";
            when "1111110101" => data <= "01110111010111011000";
            when "1111110110" => data <= "01111000000111100100";
            when "1111110111" => data <= "01111000110111110010";
            when "1111111000" => data <= "01111001100111111111";
            when "1111111001" => data <= "01111010101000001101";
            when "1111111010" => data <= "01111011011000011010";
            when "1111111011" => data <= "01111100001000100110";
            when "1111111100" => data <= "01111100111000110001";
            when "1111111101" => data <= "01111101101000111001";
            when "1111111110" => data <= "01111110011001000000";
            when others       => data <= "01111111001001000100";
        end case;
    end process rom;

end platform_independent;